parameter BUFFER_SIZE_BITS = 11;
parameter DATA_WIDTH_BITS = 16;
parameter MAX_TAU = 40;
parameter THRESHOLD = 1;
parameter WINDOW_SIZE_BITS = 8; // W = 256 